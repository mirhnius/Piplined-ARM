module InstructionMeM(input [31:0]  PC, output reg [31:0] Instruction);
  always @(PC) begin
    case (PC)
      0: Instruction <= 32'b11100011101000000000000000010100;
      4: Instruction <= 32'b11100011101000000001101000000001;
      8: Instruction <= 32'b11100011101000000010000100000011;
      12: Instruction <= 32'b11100000100100100011000000000010;
      16: Instruction <= 32'b11100000101000000100000000000000;
      20: Instruction <= 32'b11100000010001000101000100000100;
      24: Instruction <= 32'b11100000110000000110000010100000;
      28: Instruction <= 32'b11100001100001010111000101000010;
      32: Instruction <= 32'b11100000000001111000000000000011;
      36: Instruction <= 32'b11100001111000001001000000000110;
      40: Instruction <= 32'b11100000001001001010000000000101;
      44: Instruction <= 32'b11100001010110000000000000000110;
      48: Instruction <= 32'b00010000100000010001000000000001;
      52: Instruction <= 32'b11100001000110010000000000001000;
      56: Instruction <= 32'b00000000100000100010000000000010;
      60: Instruction <= 32'b11100011101000000000101100000001;
      64: Instruction <= 32'b11100100100000000001000000000000;
      68: Instruction <= 32'b11100100100100001011000000000000;
      72: Instruction <= 32'b11100100100000000010000000000100;
      76: Instruction <= 32'b11100100100000000011000000001000;
      80: Instruction <= 32'b11100100100000000100000000001101;
      84: Instruction <= 32'b11100100100000000101000000010000;
      88: Instruction <= 32'b11100100100000000110000000010100;
      92: Instruction <= 32'b11100100100100001010000000000100;
      96: Instruction <= 32'b11100100100000000111000000011000;
      100: Instruction <= 32'b11100011101000000001000000000100;
      104: Instruction <= 32'b11100011101000000010000000000000;
      108: Instruction <= 32'b11100011101000000011000000000000;
      112: Instruction <= 32'b11100000100000000100000100000011;
      116: Instruction <= 32'b11100100100101000101000000000000;
      120: Instruction <= 32'b11100100100101000110000000000100;
      124: Instruction <= 32'b11100001010101010000000000000110;
      128: Instruction <= 32'b11000100100001000110000000000000;
      132: Instruction <= 32'b11000100100001000101000000000100;
      136: Instruction <= 32'b11100010100000110011000000000001;
      140: Instruction <= 32'b11100011010100110000000000000011;
      144: Instruction <= 32'b10111010111111111111111111110111;
      148: Instruction <= 32'b11100010100000100010000000000001;
      152: Instruction <= 32'b11100001010100100000000000000001;
      156: Instruction <= 32'b10111010111111111111111111110011;
      160: Instruction <= 32'b11100100100100000001000000000000;
      164: Instruction <= 32'b11100100100100000010000000000100;
      168: Instruction <= 32'b11100100100100000011000000001000;
      172: Instruction <= 32'b11100100100100000100000000001100;
      176: Instruction <= 32'b11100100100100000101000000010000;
      180: Instruction <= 32'b11100100100100000110000000010100;
      184: Instruction <= 32'b11101010111111111111111111111111;
      default: Instruction <= 32'b00000000000000000000000000000000;
    endcase
  end
endmodule
    
